library verilog;
use verilog.vl_types.all;
entity ID_EXE_sv_unit is
end ID_EXE_sv_unit;
